module and8 (clk, rst, Input_1, Input_2, Input_3, Input_4, Input_5, Input_6, llolkek, Input_7, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Input_1;
  input  wire [0:0] Input_2;
  input  wire [0:0] Input_3;
  input  wire [0:0] Input_4;
  input  wire [0:0] Input_5;
  input  wire [0:0] Input_6;
  input  wire [0:0] llolkek;
  input  wire [0:0] Input_7;
  output  wire [0:0] Output;

  TC_And3 # (.UUID(64'd3018018426116657090 ^ UUID), .BIT_WIDTH(64'd1)) And3_0 (.in0(wire_3), .in1(wire_6), .in2(wire_4), .out(wire_2));
  TC_And3 # (.UUID(64'd2198035730399106101 ^ UUID), .BIT_WIDTH(64'd1)) And3_1 (.in0(wire_2), .in1(wire_5), .in2(wire_9), .out(wire_10));
  TC_And3 # (.UUID(64'd3924635111503222550 ^ UUID), .BIT_WIDTH(64'd1)) And3_2 (.in0(wire_10), .in1(wire_7), .in2(wire_8), .out(wire_11));
  TC_And # (.UUID(64'd2435468719362258848 ^ UUID), .BIT_WIDTH(64'd1)) And_3 (.in0(wire_11), .in1(wire_0), .out(wire_1));

  wire [0:0] wire_0;
  assign wire_0 = llolkek;
  wire [0:0] wire_1;
  assign Output = wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  assign wire_3 = Input_7;
  wire [0:0] wire_4;
  assign wire_4 = Input_2;
  wire [0:0] wire_5;
  assign wire_5 = Input_1;
  wire [0:0] wire_6;
  assign wire_6 = Input_4;
  wire [0:0] wire_7;
  assign wire_7 = Input_5;
  wire [0:0] wire_8;
  assign wire_8 = Input_6;
  wire [0:0] wire_9;
  assign wire_9 = Input_3;
  wire [0:0] wire_10;
  wire [0:0] wire_11;

endmodule
