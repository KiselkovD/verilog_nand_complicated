module COND (clk, rst, Condition, Input, Result);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Condition;
  input  wire [7:0] Input;
  output  wire [0:0] Result;

  TC_Decoder3 # (.UUID(64'd767105559009491895 ^ UUID)) Decoder3_0 (.dis(1'd0), .sel0(wire_19), .sel1(wire_3), .sel2(wire_26), .out0(), .out1(wire_2), .out2(wire_6), .out3(wire_27), .out4(wire_15), .out5(wire_8), .out6(wire_21), .out7(wire_11));
  TC_Splitter8 # (.UUID(64'd1731687480239450725 ^ UUID)) Splitter8_1 (.in(wire_22), .out0(wire_19), .out1(wire_3), .out2(wire_26), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2763831472592138518 ^ UUID)) Splitter8_2 (.in(wire_20), .out0(wire_23), .out1(wire_5), .out2(wire_4), .out3(wire_28), .out4(wire_14), .out5(wire_0), .out6(wire_17), .out7(wire_9));
  TC_Or3 # (.UUID(64'd4238712671205480422 ^ UUID), .BIT_WIDTH(64'd1)) Or3_3 (.in0(wire_23), .in1(wire_5), .in2(wire_4), .out(wire_24));
  TC_Or3 # (.UUID(64'd1865666558648900281 ^ UUID), .BIT_WIDTH(64'd1)) Or3_4 (.in0(wire_28), .in1(wire_14), .in2(wire_0), .out(wire_29));
  TC_Or # (.UUID(64'd122134950752033172 ^ UUID), .BIT_WIDTH(64'd1)) Or_5 (.in0(wire_17), .in1(wire_9), .out(wire_12));
  TC_Or3 # (.UUID(64'd2540803238069716805 ^ UUID), .BIT_WIDTH(64'd1)) Or3_6 (.in0(wire_24), .in1(wire_29), .in2(wire_12), .out(wire_16));
  TC_Not # (.UUID(64'd2066720155740043421 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_16), .out(wire_18));
  TC_Switch # (.UUID(64'd1645427440068343036 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_8 (.en(wire_6), .in(wire_9), .out(wire_7_4));
  TC_Switch # (.UUID(64'd2331709893331206764 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_9 (.en(wire_27), .in(wire_13), .out(wire_7_3));
  TC_Switch # (.UUID(64'd2338246113426213500 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_10 (.en(wire_15), .in(wire_10), .out(wire_7_5));
  TC_Switch # (.UUID(64'd1673698140392567740 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_8), .in(wire_16), .out(wire_7_0));
  TC_Switch # (.UUID(64'd2001400884787593023 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_12 (.en(wire_21), .in(wire_25), .out(wire_7_6));
  TC_Switch # (.UUID(64'd3249154913394797867 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_13 (.en(wire_11), .in(wire_1), .out(wire_7_2));
  TC_Switch # (.UUID(64'd580625633399087524 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_2), .in(wire_18), .out(wire_7_1));
  TC_Not # (.UUID(64'd3400530365242311311 ^ UUID), .BIT_WIDTH(64'd1)) Not_15 (.in(wire_9), .out(wire_25));
  TC_Not # (.UUID(64'd4066677469029232307 ^ UUID), .BIT_WIDTH(64'd1)) Not_16 (.in(wire_13), .out(wire_1));
  TC_Constant # (.UUID(64'd1318776730740804378 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out(wire_10));
  TC_Or # (.UUID(64'd2290584802158228835 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_18), .in1(wire_9), .out(wire_13));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_7_0;
  wire [0:0] wire_7_1;
  wire [0:0] wire_7_2;
  wire [0:0] wire_7_3;
  wire [0:0] wire_7_4;
  wire [0:0] wire_7_5;
  wire [0:0] wire_7_6;
  assign wire_7 = wire_7_0|wire_7_1|wire_7_2|wire_7_3|wire_7_4|wire_7_5|wire_7_6;
  assign Result = wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  assign wire_20 = Input;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  assign wire_22 = Condition;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;

endmodule
