module CPU (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input;
  output  wire [7:0] Output;

  TC_Decoder3 # (.UUID(64'd789462161731707770 ^ UUID)) Decoder3_0 (.dis(wire_10), .sel0(wire_38), .sel1(wire_34), .sel2(wire_23), .out0(wire_30), .out1(wire_4), .out2(wire_6), .out3(wire_3), .out4(wire_28), .out5(wire_20), .out6(wire_12), .out7());
  TC_Decoder3 # (.UUID(64'd2463885457538766482 ^ UUID)) Decoder3_1 (.dis(wire_10), .sel0(wire_14), .sel1(wire_33), .sel2(wire_5), .out0(wire_37), .out1(wire_18), .out2(wire_11), .out3(wire_35), .out4(wire_22), .out5(wire_31), .out6(wire_0), .out7());
  TC_Splitter8 # (.UUID(64'd4127507573354610641 ^ UUID)) Splitter8_2 (.in(wire_1), .out0(wire_38), .out1(wire_34), .out2(wire_23), .out3(wire_14), .out4(wire_33), .out5(wire_5), .out6(), .out7());
  TC_Not # (.UUID(64'd4016597418867286406 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_32), .out(wire_10));
  TC_Or # (.UUID(64'd3471351627487651955 ^ UUID), .BIT_WIDTH(64'd1)) Or_4 (.in0(wire_3), .in1(wire_7), .out(wire_21));
  TC_Mux # (.UUID(64'd1866316232879883734 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_5 (.sel(wire_7), .in0(wire_2), .in1(wire_8), .out(wire_26));
  TC_Counter # (.UUID(64'd919271322122277429 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_6 (.clk(clk), .rst(rst), .save(wire_25), .in(wire_36), .out(wire_16));
  TC_Or # (.UUID(64'd1934878915714558152 ^ UUID), .BIT_WIDTH(64'd1)) Or_7 (.in0(wire_30), .in1(wire_13), .out(wire_15));
  TC_Mux # (.UUID(64'd2860512883322327249 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_8 (.sel(wire_13), .in0(wire_2), .in1(wire_1), .out(wire_19));
  TC_And # (.UUID(64'd330084912507501615 ^ UUID), .BIT_WIDTH(64'd1)) And_9 (.in0(wire_29), .in1(wire_27), .out(wire_25));
  TC_Switch # (.UUID(64'd2775582871351875648 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_10 (.en(wire_12), .in(wire_2), .out(Output));
  TC_Switch # (.UUID(64'd4044376122156023687 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_0), .in(wire_39), .out(wire_2_6));
  DEC # (.UUID(64'd2459609941860001208 ^ UUID)) DEC_12 (.clk(clk), .rst(rst), .OPCODE(wire_1), .IMMEDIATE(wire_13), .CALCULATION(wire_7), .COPY(wire_32), .CONDITION(wire_27));
  ALU # (.UUID(64'd17775550716235650 ^ UUID)) ALU_13 (.clk(clk), .rst(rst), .Instruction(wire_1), .Input_1(wire_17), .Input_2(wire_9), .Output(wire_8));
  RegisterPlus # (.UUID(64'd156112890976078798 ^ UUID)) RegisterPlus_14 (.clk(clk), .rst(rst), .Load(wire_37), .Save_value(wire_19), .Save(wire_15), .Always_output(wire_36), .Output(wire_2_2));
  RegisterPlus # (.UUID(64'd4464545246616181500 ^ UUID)) RegisterPlus_15 (.clk(clk), .rst(rst), .Load(wire_18), .Save_value(wire_2), .Save(wire_4), .Always_output(wire_17), .Output(wire_2_5));
  RegisterPlus # (.UUID(64'd3930106220575007809 ^ UUID)) RegisterPlus_16 (.clk(clk), .rst(rst), .Load(wire_11), .Save_value(wire_2), .Save(wire_6), .Always_output(wire_9), .Output(wire_2_3));
  RegisterPlus # (.UUID(64'd552432858237882774 ^ UUID)) RegisterPlus_17 (.clk(clk), .rst(rst), .Load(wire_35), .Save_value(wire_26), .Save(wire_21), .Always_output(wire_24), .Output(wire_2_1));
  RegisterPlus # (.UUID(64'd4308030715466344996 ^ UUID)) RegisterPlus_18 (.clk(clk), .rst(rst), .Load(wire_22), .Save_value(wire_2), .Save(wire_28), .Always_output(), .Output(wire_2_4));
  RegisterPlus # (.UUID(64'd87567289778655056 ^ UUID)) RegisterPlus_19 (.clk(clk), .rst(rst), .Load(wire_31), .Save_value(wire_2), .Save(wire_20), .Always_output(), .Output(wire_2_0));
  COND_2 # (.UUID(64'd1536425055328680480 ^ UUID)) COND_2_20 (.clk(clk), .rst(rst), .Condition(wire_1), .Input(wire_24), .Result(wire_29));
  PROG # (.UUID(64'd1197309301388125823 ^ UUID)) PROG_21 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_1));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  wire [7:0] wire_2_6;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [7:0] wire_39;
  assign wire_39 = Input;

endmodule
