module ALU (clk, rst, Instruction, Input_1, Input_2, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Instruction;
  input  wire [7:0] Input_1;
  input  wire [7:0] Input_2;
  output  wire [7:0] Output;

  TC_Splitter8 # (.UUID(64'd4321707480502513143 ^ UUID)) Splitter8_0 (.in(wire_23), .out0(wire_11), .out1(wire_7), .out2(wire_25), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd1047726087564551862 ^ UUID)) Decoder3_1 (.dis(1'd0), .sel0(wire_11), .sel1(wire_7), .sel2(wire_25), .out0(wire_2), .out1(wire_20), .out2(wire_10), .out3(wire_19), .out4(wire_9), .out5(wire_21), .out6(), .out7());
  TC_Or # (.UUID(64'd3697877361305982650 ^ UUID), .BIT_WIDTH(64'd8)) Or8_2 (.in0(wire_3), .in1(wire_6), .out(wire_12));
  TC_Not # (.UUID(64'd2017182251518901485 ^ UUID), .BIT_WIDTH(64'd8)) Not8_3 (.in(wire_6), .out(wire_15));
  TC_Or # (.UUID(64'd3579128892170319245 ^ UUID), .BIT_WIDTH(64'd8)) Or8_4 (.in0(wire_22), .in1(wire_15), .out(wire_0));
  TC_Switch # (.UUID(64'd1838319591841633892 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_2), .in(wire_12), .out(wire_4_0));
  TC_Switch # (.UUID(64'd2254496928853479681 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_10), .in(wire_14), .out(wire_4_2));
  TC_Switch # (.UUID(64'd396306721349376195 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_19), .in(wire_1), .out(wire_4_3));
  TC_Switch # (.UUID(64'd4538812189126161630 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_20), .in(wire_0), .out(wire_4_5));
  TC_Not # (.UUID(64'd1286176436029887504 ^ UUID), .BIT_WIDTH(64'd8)) Not8_9 (.in(wire_3), .out(wire_22));
  TC_Not # (.UUID(64'd1738053492834767768 ^ UUID), .BIT_WIDTH(64'd8)) Not8_10 (.in(wire_16), .out(wire_14));
  TC_Not # (.UUID(64'd287793528915418250 ^ UUID), .BIT_WIDTH(64'd8)) Not8_11 (.in(wire_3), .out(wire_13));
  TC_Not # (.UUID(64'd1166442119747664101 ^ UUID), .BIT_WIDTH(64'd8)) Not8_12 (.in(wire_6), .out(wire_5));
  TC_Or # (.UUID(64'd1842676259106870302 ^ UUID), .BIT_WIDTH(64'd8)) Or8_13 (.in0(wire_3), .in1(wire_6), .out(wire_16));
  TC_Not # (.UUID(64'd389128709749653788 ^ UUID), .BIT_WIDTH(64'd8)) Not8_14 (.in(wire_17), .out(wire_1));
  TC_Or # (.UUID(64'd638383184506304288 ^ UUID), .BIT_WIDTH(64'd8)) Or8_15 (.in0(wire_13), .in1(wire_5), .out(wire_17));
  TC_Switch # (.UUID(64'd4541383247443122317 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_9), .in(wire_24), .out(wire_4_1));
  TC_Switch # (.UUID(64'd4225945799929144992 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_21), .in(wire_8), .out(wire_4_4));
  TC_Add # (.UUID(64'd2623997479491979901 ^ UUID), .BIT_WIDTH(64'd8)) Add8_18 (.in0(wire_3), .in1(wire_6), .ci(1'd0), .out(wire_24), .co());
  TC_Add # (.UUID(64'd2415820346936528038 ^ UUID), .BIT_WIDTH(64'd8)) Add8_19 (.in0(wire_3), .in1(wire_18), .ci(1'd0), .out(wire_8), .co());
  TC_Neg # (.UUID(64'd2828099826108676478 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_20 (.in(wire_6), .out(wire_18));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  assign wire_3 = Input_1;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  wire [7:0] wire_4_4;
  wire [7:0] wire_4_5;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5;
  assign Output = wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  assign wire_6 = Input_2;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_23;
  assign wire_23 = Instruction;
  wire [7:0] wire_24;
  wire [0:0] wire_25;

endmodule
