module PROG (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input;
  output  wire [7:0] Output;

  TC_Splitter8 # (.UUID(64'd2435112095298298361 ^ UUID)) Splitter8_0 (.in(wire_7), .out0(wire_44), .out1(wire_31), .out2(wire_34), .out3(wire_25), .out4(), .out5(), .out6(), .out7());
  TC_Decoder1 # (.UUID(64'd2328959383735369342 ^ UUID)) Decoder1_1 (.sel(wire_44), .out0(wire_14), .out1(wire_10));
  TC_Decoder1 # (.UUID(64'd4453464714108961545 ^ UUID)) Decoder1_2 (.sel(wire_31), .out0(wire_15), .out1(wire_1));
  TC_Decoder1 # (.UUID(64'd680292653085339257 ^ UUID)) Decoder1_3 (.sel(wire_34), .out0(wire_11), .out1(wire_23));
  TC_Decoder1 # (.UUID(64'd1887189890146492707 ^ UUID)) Decoder1_4 (.sel(wire_25), .out0(wire_8), .out1(wire_12));
  RegisterPlus # (.UUID(64'd3477855810552793057 ^ UUID)) RegisterPlus_5 (.clk(clk), .rst(rst), .Load(wire_20), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_7));
  and8 # (.UUID(64'd1854568874100887990 ^ UUID)) and8_6 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_11), .Input_3(wire_13), .Input_4(wire_15), .Input_5(wire_13), .Input_6(wire_13), .llolkek(wire_13), .Input_7(wire_14), .Output(wire_20));
  TC_Constant # (.UUID(64'd2568444835643953338 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out(wire_13));
  RegisterPlus # (.UUID(64'd55276178600414620 ^ UUID)) RegisterPlus_8 (.clk(clk), .rst(rst), .Load(wire_42), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_4));
  and8 # (.UUID(64'd1961325811558144586 ^ UUID)) and8_9 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_11), .Input_3(wire_26), .Input_4(wire_15), .Input_5(wire_26), .Input_6(wire_26), .llolkek(wire_26), .Input_7(wire_10), .Output(wire_42));
  TC_Constant # (.UUID(64'd421430877386728711 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out(wire_26));
  RegisterPlus # (.UUID(64'd2863992784825382537 ^ UUID)) RegisterPlus_11 (.clk(clk), .rst(rst), .Load(wire_30), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_5));
  and8 # (.UUID(64'd736316101638821330 ^ UUID)) and8_12 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_11), .Input_3(wire_43), .Input_4(wire_1), .Input_5(wire_43), .Input_6(wire_43), .llolkek(wire_43), .Input_7(wire_14), .Output(wire_30));
  TC_Constant # (.UUID(64'd2632105423500060957 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out(wire_43));
  RegisterPlus # (.UUID(64'd3152801442508544873 ^ UUID)) RegisterPlus_14 (.clk(clk), .rst(rst), .Load(wire_27), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_13));
  and8 # (.UUID(64'd559851590864566962 ^ UUID)) and8_15 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_11), .Input_3(wire_22), .Input_4(wire_1), .Input_5(wire_22), .Input_6(wire_22), .llolkek(wire_22), .Input_7(wire_10), .Output(wire_27));
  TC_Constant # (.UUID(64'd1632033517224195888 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_22));
  RegisterPlus # (.UUID(64'd686901985730980529 ^ UUID)) RegisterPlus_17 (.clk(clk), .rst(rst), .Load(wire_41), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_2));
  and8 # (.UUID(64'd2038290010876050318 ^ UUID)) and8_18 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_23), .Input_3(wire_5), .Input_4(wire_15), .Input_5(wire_5), .Input_6(wire_5), .llolkek(wire_5), .Input_7(wire_14), .Output(wire_41));
  TC_Constant # (.UUID(64'd1319027891604423226 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_19 (.out(wire_5));
  RegisterPlus # (.UUID(64'd3001945359049208787 ^ UUID)) RegisterPlus_20 (.clk(clk), .rst(rst), .Load(wire_45), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_6));
  and8 # (.UUID(64'd1690636845594045670 ^ UUID)) and8_21 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_23), .Input_3(wire_9), .Input_4(wire_15), .Input_5(wire_9), .Input_6(wire_9), .llolkek(wire_9), .Input_7(wire_10), .Output(wire_45));
  TC_Constant # (.UUID(64'd2889423854709821689 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_22 (.out(wire_9));
  RegisterPlus # (.UUID(64'd495269329642429205 ^ UUID)) RegisterPlus_23 (.clk(clk), .rst(rst), .Load(wire_37), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_11));
  and8 # (.UUID(64'd2327651323208194487 ^ UUID)) and8_24 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_23), .Input_3(wire_6), .Input_4(wire_1), .Input_5(wire_6), .Input_6(wire_6), .llolkek(wire_6), .Input_7(wire_14), .Output(wire_37));
  TC_Constant # (.UUID(64'd4356675971236521367 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out(wire_6));
  RegisterPlus # (.UUID(64'd1545498608926041819 ^ UUID)) RegisterPlus_26 (.clk(clk), .rst(rst), .Load(wire_28), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_9));
  and8 # (.UUID(64'd3633203500260515148 ^ UUID)) and8_27 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_23), .Input_3(wire_0), .Input_4(wire_1), .Input_5(wire_0), .Input_6(wire_0), .llolkek(wire_0), .Input_7(wire_10), .Output(wire_28));
  TC_Constant # (.UUID(64'd2410756799956088170 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_28 (.out(wire_0));
  RegisterPlus # (.UUID(64'd1739888728747161338 ^ UUID)) RegisterPlus_29 (.clk(clk), .rst(rst), .Load(wire_39), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_15));
  and8 # (.UUID(64'd3260625674356521876 ^ UUID)) and8_30 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_11), .Input_3(wire_4), .Input_4(wire_15), .Input_5(wire_4), .Input_6(wire_4), .llolkek(wire_4), .Input_7(wire_10), .Output(wire_39));
  TC_Constant # (.UUID(64'd4317447753839421711 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_31 (.out(wire_4));
  RegisterPlus # (.UUID(64'd796689678003878509 ^ UUID)) RegisterPlus_32 (.clk(clk), .rst(rst), .Load(wire_36), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_3));
  and8 # (.UUID(64'd1129499025503222550 ^ UUID)) and8_33 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_11), .Input_3(wire_35), .Input_4(wire_1), .Input_5(wire_35), .Input_6(wire_35), .llolkek(wire_35), .Input_7(wire_14), .Output(wire_36));
  TC_Constant # (.UUID(64'd969447812076161726 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_34 (.out(wire_35));
  RegisterPlus # (.UUID(64'd758671467874901218 ^ UUID)) RegisterPlus_35 (.clk(clk), .rst(rst), .Load(wire_17), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_0));
  and8 # (.UUID(64'd3796142071410602525 ^ UUID)) and8_36 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_11), .Input_3(wire_24), .Input_4(wire_1), .Input_5(wire_24), .Input_6(wire_24), .llolkek(wire_24), .Input_7(wire_10), .Output(wire_17));
  TC_Constant # (.UUID(64'd36991073773931435 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_37 (.out(wire_24));
  RegisterPlus # (.UUID(64'd2600144778229742400 ^ UUID)) RegisterPlus_38 (.clk(clk), .rst(rst), .Load(wire_40), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_8));
  and8 # (.UUID(64'd2092619706795044061 ^ UUID)) and8_39 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_23), .Input_3(wire_18), .Input_4(wire_15), .Input_5(wire_18), .Input_6(wire_18), .llolkek(wire_18), .Input_7(wire_14), .Output(wire_40));
  TC_Constant # (.UUID(64'd1239211769493268583 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_40 (.out(wire_18));
  RegisterPlus # (.UUID(64'd3540119006208166081 ^ UUID)) RegisterPlus_41 (.clk(clk), .rst(rst), .Load(wire_21), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_14));
  and8 # (.UUID(64'd1979992577759958344 ^ UUID)) and8_42 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_23), .Input_3(wire_2), .Input_4(wire_15), .Input_5(wire_2), .Input_6(wire_2), .llolkek(wire_2), .Input_7(wire_10), .Output(wire_21));
  TC_Constant # (.UUID(64'd148066942694921782 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_43 (.out(wire_2));
  RegisterPlus # (.UUID(64'd1188714155507598778 ^ UUID)) RegisterPlus_44 (.clk(clk), .rst(rst), .Load(wire_32), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_1));
  and8 # (.UUID(64'd4362869593957121707 ^ UUID)) and8_45 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_23), .Input_3(wire_29), .Input_4(wire_1), .Input_5(wire_29), .Input_6(wire_29), .llolkek(wire_29), .Input_7(wire_14), .Output(wire_32));
  TC_Constant # (.UUID(64'd1836366440658814316 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_46 (.out(wire_29));
  RegisterPlus # (.UUID(64'd4259648734336962092 ^ UUID)) RegisterPlus_47 (.clk(clk), .rst(rst), .Load(wire_38), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_10));
  and8 # (.UUID(64'd1512921030119820249 ^ UUID)) and8_48 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_23), .Input_3(wire_19), .Input_4(wire_1), .Input_5(wire_19), .Input_6(wire_19), .llolkek(wire_19), .Input_7(wire_10), .Output(wire_38));
  TC_Constant # (.UUID(64'd370263691251949185 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_49 (.out(wire_19));
  RegisterPlus # (.UUID(64'd4117960188568936424 ^ UUID)) RegisterPlus_50 (.clk(clk), .rst(rst), .Load(wire_33), .Save_value(8'd0), .Save(1'd0), .Always_output(), .Output(wire_3_12));
  and8 # (.UUID(64'd256384586740577307 ^ UUID)) and8_51 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_11), .Input_3(wire_16), .Input_4(wire_15), .Input_5(wire_16), .Input_6(wire_16), .llolkek(wire_16), .Input_7(wire_14), .Output(wire_33));
  TC_Constant # (.UUID(64'd3920281642702204061 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_52 (.out(wire_16));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  wire [7:0] wire_3_8;
  wire [7:0] wire_3_9;
  wire [7:0] wire_3_10;
  wire [7:0] wire_3_11;
  wire [7:0] wire_3_12;
  wire [7:0] wire_3_13;
  wire [7:0] wire_3_14;
  wire [7:0] wire_3_15;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7|wire_3_8|wire_3_9|wire_3_10|wire_3_11|wire_3_12|wire_3_13|wire_3_14|wire_3_15;
  assign Output = wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = Input;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;

endmodule
